  --Example instantiation for system 'unnamed'
  unnamed_inst : unnamed
    port map(
      out_pwm_from_the_avalon_pwm_0 => out_pwm_from_the_avalon_pwm_0,
      clk_0 => clk_0,
      reset_n => reset_n
    );


